module o_logic();
    input	[1:0]	gp1;
	input	[1:0]	gp2;
	output	[1:0]	r;


endmodule