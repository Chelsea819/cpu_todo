/*************************************************************************
	> File Name: add.v
	> Author: Chelsea
	> Mail: 1938166340@qq.com 
	> Created Time: 2024年04月16日 星期二 15时59分48秒
 ************************************************************************/

module ysyx_22041211_ (
);


